module val

pub interface Struct {
}
