module val

pub type Uint = u8 | u16 | u32 | u64
