module val

pub type Int = byte
	| u16
	| u32
	| u64
	| i8
	| i16
	| int // alias i32
	| i64
