module val

pub type Float = f32 | f64
