module val

pub struct Nil {}

pub interface Struct {
}
