module val

pub type Number = byte | u16 | u32 | u64 | i8 | i16 | int | i64 | f32 | f64
