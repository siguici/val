module val

pub type Uint = byte // alias u8
	| u16
	| u32
	| u64
