module val

import time

pub type Primitive = Nil
	| voidptr
	| bool
	| byte
	| u16
	| u32
	| u64
	| i8
	| i16
	| int
	| i64
	| f32
	| f64
	| rune
	| string
	| time.Time
	| []Primitive
